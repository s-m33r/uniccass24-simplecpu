magic
tech sky130A
magscale 1 2
timestamp 1729498058
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 76 558808 349840
<< metal2 >>
rect 19154 0 19210 800
rect 56414 0 56470 800
rect 93674 0 93730 800
rect 130934 0 130990 800
rect 168194 0 168250 800
rect 205454 0 205510 800
rect 242714 0 242770 800
rect 279974 0 280030 800
rect 317234 0 317290 800
rect 354494 0 354550 800
rect 391754 0 391810 800
rect 429014 0 429070 800
rect 466274 0 466330 800
rect 503534 0 503590 800
rect 540794 0 540850 800
<< obsm2 >>
rect 4214 856 558514 349829
rect 4214 70 19098 856
rect 19266 70 56358 856
rect 56526 70 93618 856
rect 93786 70 130878 856
rect 131046 70 168138 856
rect 168306 70 205398 856
rect 205566 70 242658 856
rect 242826 70 279918 856
rect 280086 70 317178 856
rect 317346 70 354438 856
rect 354606 70 391698 856
rect 391866 70 428958 856
rect 429126 70 466218 856
rect 466386 70 503478 856
rect 503646 70 540738 856
rect 540906 70 558514 856
<< metal3 >>
rect 559200 338920 560000 339040
rect 559200 317160 560000 317280
rect 559200 295400 560000 295520
rect 559200 273640 560000 273760
rect 559200 251880 560000 252000
rect 559200 230120 560000 230240
rect 559200 208360 560000 208480
rect 559200 186600 560000 186720
rect 559200 164840 560000 164960
rect 559200 143080 560000 143200
rect 559200 121320 560000 121440
rect 559200 99560 560000 99680
rect 559200 77800 560000 77920
rect 559200 56040 560000 56160
rect 559200 34280 560000 34400
rect 559200 12520 560000 12640
<< obsm3 >>
rect 4210 339120 559200 349825
rect 4210 338840 559120 339120
rect 4210 317360 559200 338840
rect 4210 317080 559120 317360
rect 4210 295600 559200 317080
rect 4210 295320 559120 295600
rect 4210 273840 559200 295320
rect 4210 273560 559120 273840
rect 4210 252080 559200 273560
rect 4210 251800 559120 252080
rect 4210 230320 559200 251800
rect 4210 230040 559120 230320
rect 4210 208560 559200 230040
rect 4210 208280 559120 208560
rect 4210 186800 559200 208280
rect 4210 186520 559120 186800
rect 4210 165040 559200 186520
rect 4210 164760 559120 165040
rect 4210 143280 559200 164760
rect 4210 143000 559120 143280
rect 4210 121520 559200 143000
rect 4210 121240 559120 121520
rect 4210 99760 559200 121240
rect 4210 99480 559120 99760
rect 4210 78000 559200 99480
rect 4210 77720 559120 78000
rect 4210 56240 559200 77720
rect 4210 55960 559120 56240
rect 4210 34480 559200 55960
rect 4210 34200 559120 34480
rect 4210 12720 559200 34200
rect 4210 12440 559120 12720
rect 4210 1259 559200 12440
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 449387 2048 449568 15333
rect 450048 2048 464928 15333
rect 465408 2048 479445 15333
rect 449387 1939 479445 2048
<< labels >>
rlabel metal3 s 559200 34280 560000 34400 6 io_oeb[0]
port 1 nsew signal output
rlabel metal3 s 559200 77800 560000 77920 6 io_oeb[1]
port 2 nsew signal output
rlabel metal3 s 559200 121320 560000 121440 6 io_oeb[2]
port 3 nsew signal output
rlabel metal3 s 559200 164840 560000 164960 6 io_oeb[3]
port 4 nsew signal output
rlabel metal3 s 559200 208360 560000 208480 6 io_oeb[4]
port 5 nsew signal output
rlabel metal3 s 559200 251880 560000 252000 6 io_oeb[5]
port 6 nsew signal output
rlabel metal3 s 559200 295400 560000 295520 6 io_oeb[6]
port 7 nsew signal output
rlabel metal3 s 559200 338920 560000 339040 6 io_oeb[7]
port 8 nsew signal output
rlabel metal3 s 559200 12520 560000 12640 6 io_out[0]
port 9 nsew signal output
rlabel metal3 s 559200 56040 560000 56160 6 io_out[1]
port 10 nsew signal output
rlabel metal3 s 559200 99560 560000 99680 6 io_out[2]
port 11 nsew signal output
rlabel metal3 s 559200 143080 560000 143200 6 io_out[3]
port 12 nsew signal output
rlabel metal3 s 559200 186600 560000 186720 6 io_out[4]
port 13 nsew signal output
rlabel metal3 s 559200 230120 560000 230240 6 io_out[5]
port 14 nsew signal output
rlabel metal3 s 559200 273640 560000 273760 6 io_out[6]
port 15 nsew signal output
rlabel metal3 s 559200 317160 560000 317280 6 io_out[7]
port 16 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_in[0]
port 17 nsew signal input
rlabel metal2 s 429014 0 429070 800 6 la_data_in[10]
port 18 nsew signal input
rlabel metal2 s 466274 0 466330 800 6 la_data_in[11]
port 19 nsew signal input
rlabel metal2 s 503534 0 503590 800 6 la_data_in[12]
port 20 nsew signal input
rlabel metal2 s 540794 0 540850 800 6 la_data_in[13]
port 21 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[1]
port 22 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_data_in[3]
port 24 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_data_in[4]
port 25 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_data_in[5]
port 26 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_data_in[6]
port 27 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_data_in[7]
port 28 nsew signal input
rlabel metal2 s 354494 0 354550 800 6 la_data_in[8]
port 29 nsew signal input
rlabel metal2 s 391754 0 391810 800 6 la_data_in[9]
port 30 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 32 nsew ground bidirectional
rlabel metal2 s 19154 0 19210 800 6 wb_clk_i
port 33 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 55096798
string GDS_FILE /home/labuser/uniccass24-simplecpu/openlane/user_proj_example/runs/24_10_21_13_29/results/signoff/user_proj_example.magic.gds
string GDS_START 594808
<< end >>

